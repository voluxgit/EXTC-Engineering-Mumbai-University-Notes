*** SPICE deck for cell expt2{sch} from library expt2
*** Created on Sun Nov 06, 2022 17:33:47
*** Last revised on Sun Nov 06, 2022 18:19:24
*** Written on Sun Nov 06, 2022 20:08:12 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: expt2{sch}
Mnmos@0 out in gnd gnd NMOS L=0.6U W=3U
Mpmos@0 vdd in out vdd PMOS L=0.6U W=3U

* Spice Code nodes in cell cell 'expt2{sch}'
vdd vdd 0 DC 5
vin in 0 DC pwl 10n 0 20n 5 50n 5 60n 0
cload out 0 250fF
.measure tran tf trig v(out) val=4.5 fall=1 td=8ns targ v(out) val=0.5 fall=1
.measure tran tr trig v(out) val=0.5 rise=1 td=50ns targ v(out) val=4.5 rise=1
.tran 0 100ns
.include D:\college related\Third year\electric main\C5_models.txt
.END
